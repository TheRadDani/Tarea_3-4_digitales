module and_gate(input A, input B, output out_and_gate);
    assign #(1:2:3,1:2:3) 
    out_and_gate = A & B;
endmodule
//precio 0.90$