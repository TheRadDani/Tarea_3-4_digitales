module and_gate(output out_and_gate, input A, input B);
    assign #(1:2:3,1:2:3) out_and_gate = A & B;
endmodule
//precio 0.90$