module and_gate(output reg out_and_gate, input A, input B);
    assign #(3.5:3.5:5.9,3.5:3.5:5.9) 
    and(out_and_gate,A,B);
endmodule
//precio 0.90$